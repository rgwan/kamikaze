/* 写回寄存器与访存 */
module kamikaze_writeback(clk_i,
			rst_i);
	input clk_i;
	input rst_i;
	
	
endmodule
