module kamikaze_execute(clk_i,
			rst_i);
	input clk_i;
	input rst_i;
endmodule
